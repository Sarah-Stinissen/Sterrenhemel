library IEEE;						-- Bibliotheek ingeven waar de
use IEEE.std_logic_1164.all;		-- VHDL codes zich bevinden.
use IEEE.std_logic_unsigned.all;

entity decoder is						-- Beschrijving van schakeling.
	port(								-- In en uitgangen weergeven.
        	code_in: 	in std_logic_vector (5 downto 0);	-- 6-bits code
			code_uit:	out std_logic_vector (63 downto 0)	-- 64- bits code
		);
end decoder;								-- Einde beschrijving.

architecture gedrag of decoder is			-- Beschrijving van hardware.
begin										-- Begin hardware beschrijving.
  process(code_in)							-- Process van 6-bits naar 64-bits omvormer.
  begin										-- Begin van hardware beschrijving
    case code_in is
      	when "011000" => code_uit <=	"1111111111111111111111111111111111111111111111111111111111111110";		-- Uitgang 1  
      	when "100000" => code_uit <=	"1111111111111111111111111111111111111111111111111111111111111101";		-- Uitgang 2   
		when "110000" => code_uit <= 	"1111111111111111111111111111111111111111111111111111111111111011"; 	-- Uitgang 3  
      	when "001001" => code_uit <= 	"1111111111111111111111111111111111111111111111111111111111110111";		-- Uitgang 4  
		when "110001" => code_uit <=	"1111111111111111111111111111111111111111111111111111111111101111";		-- Uitgang 5   
		when "000110" => code_uit <= 	"1111111111111111111111111111111111111111111111111111111111011111";		-- Uitgang 6  
		when "000000" => code_uit <= 	"1111111111111111111111111111111111111111111111111111111110111111";		-- Uitgang 7   
		when "001110" => code_uit <= 	"1111111111111111111111111111111111111111111111111111111101111111";		-- Uitgang 8   
		when "001011" => code_uit <= 	"1111111111111111111111111111111111111111111111111111111011111111";		-- Uitgang 9   
		when "000001" => code_uit <= 	"1111111111111111111111111111111111111111111111111111110111111111";		-- Uitgang 10   
		when "101011" => code_uit <= 	"1111111111111111111111111111111111111111111111111111101111111111";		-- Uitgang 11 
		when "110100" => code_uit <= 	"1111111111111111111111111111111111111111111111111111011111111111";		-- Uitgang 12 
		when "001101" => code_uit <=	"1111111111111111111111111111111111111111111111111110111111111111";		-- Uitgang 13 
		when "010101" => code_uit <= 	"1111111111111111111111111111111111111111111111111101111111111111";		-- Uitgang 14 
		when "101001" => code_uit <= 	"1111111111111111111111111111111111111111111111110111111111111111";		-- Uitgang 16 
		when "010010" => code_uit <= 	"1111111111111111111111111111111111111111111111101111111111111111";		-- Uitgang 17 
		when "100010" => code_uit <=	"1111111111111111111111111111111111111111111111011111111111111111";		-- Uitgang 18 
		when "100011" => code_uit <= 	"1111111111111111111111111111111111111111111110111111111111111111";		-- Uitgang 19  
		when "011101" => code_uit <= 	"1111111111111111111111111111111111111111111101111111111111111111";		-- Uitgang 20   
		when "100101" => code_uit <= 	"1111111111111111111111111111111111111111111011111111111111111111";		-- Uitgang 21 
		when "000011" => code_uit <= 	"1111111111111111111111111111111111111111110111111111111111111111";		-- Uitgang 22 
		when "101010" => code_uit <=  	"1111111111111111111111111111111111111111101111111111111111111111";		-- Uitgang 23 
		when "001100" => code_uit <=  	"1111111111111111111111111111111111111111011111111111111111111111";		-- Uitgang 24 
		when "010011" => code_uit <= 	"1111111111111111111111111111111111111110111111111111111111111111";		-- Uitgang 25  
		when "010110" => code_uit <=  	"1111111111111111111111111111111111111101111111111111111111111111";		-- Uitgang 26 
		when "000101" => code_uit <= 	"1111111111111111111111111111111111111011111111111111111111111111";		-- Uitgang 27  
		when "100100" => code_uit <=  	"1111111111111111111111111111111111110111111111111111111111111111";		-- Uitgang 28 
		when "101110" => code_uit <=  	"1111111111111111111111111111111111101111111111111111111111111111";		-- Uitgang 29 
		when "110010" => code_uit <= 	"1111111111111111111111111111111111011111111111111111111111111111";		-- Uitgang 30  
		when "011110" => code_uit <=  	"1111111111111111111111111111111110111111111111111111111111111111";		-- Uitgang 31 
		when "011001" => code_uit <= 	"1111111111111111111111111111111101111111111111111111111111111111";		-- Uitgang 32  
		when "110011" => code_uit <=  	"1111111111111111111111111111111011111111111111111111111111111111";		-- Uitgang 33 
		when "010001" => code_uit <= 	"1111111111111111111111111111110111111111111111111111111111111111";		-- Uitgang 34  
		when "000010" => code_uit <=  	"1111111111111111111111111111101111111111111111111111111111111111";		-- Uitgang 35 
		when "101100" => code_uit <= 	"1111111111111111111111111111011111111111111111111111111111111111";		-- Uitgang 36 
		when "001010" => code_uit <=  	"1111111111111111111111111110111111111111111111111111111111111111";		-- Uitgang 37 
		when "110110" => code_uit <= 	"1111111111111111111111111101111111111111111111111111111111111111";		-- Uitgang 38  
		when "100001" => code_uit <=  	"1111111111111111111111111011111111111111111111111111111111111111";		-- Uitgang 39 
		when "100110" => code_uit <= 	"1111111111111111111111110111111111111111111111111111111111111111";		-- Uitgang 40  
		when "010100" => code_uit <=  	"1111111111111111111111101111111111111111111111111111111111111111";		-- Uitgang 41 
		when "000100" => code_uit <= 	"1111111111111111111111011111111111111111111111111111111111111111";		-- Uitgang 42  
		when "011010" => code_uit <=  	"1111111111111111111110111111111111111111111111111111111111111111";		-- Uitgang 43 
		when "101101" => code_uit <=  	"1111111111111111111101111111111111111111111111111111111111111111";		-- Uitgang 44 
		when "011011" => code_uit <= 	"1111111111111111111011111111111111111111111111111111111111111111";		-- Uitgang 45  
		when "101000" => code_uit <= 	"1111111111111111110111111111111111111111111111111111111111111111";		-- Uitgang 46  
		when "001000" => code_uit <=  	"1111111111111111101111111111111111111111111111111111111111111111";		-- Uitgang 47 
		when "010000" => code_uit <= 	"1111111111111111011111111111111111111111111111111111111111111111";		-- Uitgang 48  
		when "011100" => code_uit <=  	"1111111111111110111111111111111111111111111111111111111111111111";		-- Uitgang 49 
		when "000111" => code_uit <= 	"1111111111111101111111111111111111111111111111111111111111111111";		-- Uitgang 50  
		when "011111" => code_uit <=  	"1111111111111011111111111111111111111111111111111111111111111111";		-- Uitgang 51 
		when "001111" => code_uit <= 	"1111111111110111111111111111111111111111111111111111111111111111";		-- Uitgang 52  
		when "100111" => code_uit <=  	"1111111111101111111111111111111111111111111111111111111111111111";		-- Uitgang 53 
		when "010111" => code_uit <= 	"1111111111011111111111111111111111111111111111111111111111111111";		-- Uitgang 54  
		when "110111" => code_uit <=  	"1111111110111111111111111111111111111111111111111111111111111111";		-- Uitgang 55 
		when "101111" => code_uit <= 	"1111111101111111111111111111111111111111111111111111111111111111";		-- Uitgang 56 
		when others => code_uit <= 		"1111111111111111111111111111111111111111111111111111111111111111";		-- Anders geen enkele selecteren. 
    end case;
  end process;									-- Einde process
end;											-- Einde architecture
